module ArrayController(
    input i_clk,
    input i_rst_n,

    input i_data_valid,
    input i_dma_ready,

    output o_device_ready,
    output o_data_valid
);





endmodule